.SUBCKT C0402C102J5GACAUTO 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 10000 Hz
*KEMET Model RLC Cerm
R1 3 4 1.21294260025024
R2 2 5 0.910000026226044
R3 1 6 99999997952
L1 1 2 1.36999994682085E-11
L2 2 3 2.60299989895962E-10
C1 4 6 9.99999971718069E-10
C2 5 6 5.99999986588955E-14
.ENDS